library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Universal binary counter (ubc)
entity ubc is
   generic(N: integer := 8);
   port(
      clk, reset: in std_logic;  -- Clock and reset inputs
      en:         in std_logic;  -- Enable
      up:         in std_logic;  -- Count up or down
      max_tick, min_tick: out std_logic;
      q: out std_logic_vector(N-1 downto 0)
   );
end ubc;

architecture arch of ubc is
   signal r_reg: unsigned(N-1 downto 0);
   signal r_next: unsigned(N-1 downto 0);
begin
   -- register
   process(clk,reset)
   begin
      if (reset='1') then
         r_reg <= (others=>'0');
      elsif (clk'event and clk='1') then
         r_reg <= r_next;
      end if;
   end process;
   -- next-state logic
   r_next <= r_reg + 1     when en ='1' and up='1' else
             r_reg - 1     when en ='1' and up='0' else
             r_reg;
   -- output logic
   q <= std_logic_vector(r_reg);
   max_tick <= '1' when r_reg=(2**N-1) else '0';
   min_tick <= '1' when r_reg=0 else '0';
end arch;